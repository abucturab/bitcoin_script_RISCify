`Define OP_0 0
`Define OP_PUSHDATA1 76
`Define OP_PUSHDATA2 77
`Define OP_PUSHDATA4 78
`Define OP_1NEGATE 79
`Define OP_1 81
`Define OP_2 82
`Define OP_3 83
`Define OP_4 84
`Define OP_5 85
`Define OP_6 86
`Define OP_7 87
`Define OP_8 88
`Define OP_9 89
`Define OP_10 90
`Define OP_11 91
`Define OP_12 92
`Define OP_13 93
`Define OP_14 94
`Define OP_15 95
`Define OP_16 96
`Define OP_NOP 97
`Define OP_VER  98
`Define OP_VERIFY 105
`Define OP_RETURN 106
`Define OP_TOALTSTACK 107
`Define OP_FROMALTSTACK 108
`Define OP_2DROP 109
`Define OP_2DUP 110
`Define OP_3DUP 111
`Define OP_2OVER 112
`Define OP_2ROT 113
`Define OP_2SWAP 114
`Define OP_IFDUP 115
`Define OP_DEPTH 116
`Define OP_DROP 117
`Define OP_DUP 118
`Define OP_NIP 119
`Define OP_OVER 120
`Define OP_PICK 121
`Define OP_ROLL 122
`Define OP_ROT 123
`Define OP_SWAP 124
`Define OP_TUCK 125
`Define OP_CAT 126
`Define OP_SPLIT 127
`Define OP_NUM2BIN 128
`Define OP_BIN2NUM 129
`Define OP_SIZE 130
`Define OP_INVERT 131
`Define OP_AND 132
`Define OP_OR 133
`Define OP_XOR 134
`Define OP_EQUAL 135
`Define OP_EQUALVERIFY 136
`Define OP_1ADD 139
`Define OP_1SUB 140
`Define OP_2MUL   141
`Define OP_2DIV   142
`Define OP_NEGATE 143
`Define OP_ABS 144
`Define OP_NOT 145
`Define OP_0NOTEQUAL 146
`Define OP_ADD 147
`Define OP_SUB 148
`Define OP_MUL 149
`Define OP_DIV 150
`Define OP_MOD 151
`Define OP_LSHIFT 152
`Define OP_RSHIFT 153
`Define OP_BOOLAND 154
`Define OP_BOOLOR 155
`Define OP_NUMEQUAL 156
`Define OP_NUMEQUALVERIFY 157
`Define OP_NUMNOTEQUAL 158
`Define OP_LESSTHAN 159
`Define OP_GREATERTHAN 160
`Define OP_LESSTHANOREQUAL 161
`Define OP_GREATERTHANOREQUAL 162
`Define OP_MIN 163
`Define OP_MAX 164
`Define OP_WITHIN 165
`Define OP_RIPEMD160 166
`Define OP_SHA1 167
`Define OP_SHA256 168
`Define OP_HASH160 169
`Define OP_HASH256 170
`Define OP_CODESEPARATOR 171
`Define OP_CHECKSIG 172
`Define OP_CHECKSIGVERIFY 173
`Define OP_CHECKMULTISIG 174
`Define OP_CHECKMULTISIGVERIFY 175
`Define OP_CHECKLOCKTIMEVERIFY 177
`Define OP_CHECKSEQUENCEVERIFY 178